`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/07/2025 03:24:15 PM
// Design Name: 
// Module Name: entering_numbers
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module entering_numbers(
    input freq625m, btnC, btnU, btnL, btnR, btnD,
    output [17:0] num1, num2,
    output done);
endmodule