module font_rom(
    input [7:0] char_code,
    output reg [34:0] font_data
);

    always @(*) begin
        case (char_code)
            // Numbers
            "0": font_data = 35'b01110_10001_10011_10101_11001_10001_01110;
            "1": font_data = 35'b00100_01100_00100_00100_00100_00100_01110;
            "2": font_data = 35'b01110_10001_00001_00010_00100_01000_11111;
            "3": font_data = 35'b11111_00010_00100_00010_00001_10001_01110;
            "4": font_data = 35'b00010_00110_01010_10010_11111_00010_00010;
            "5": font_data = 35'b11111_10000_11110_00001_00001_10001_01110;
            "6": font_data = 35'b00110_01000_10000_11110_10001_10001_01110;
            "7": font_data = 35'b11111_00001_00010_00100_01000_01000_01000;
            "8": font_data = 35'b01110_10001_10001_01110_10001_10001_01110;
            "9": font_data = 35'b01110_10001_10001_01111_00001_00010_01100;
            
            // Letters
            "A": font_data = 35'b01110_10001_10001_10001_11111_10001_10001;
            "B": font_data = 35'b11110_10001_10001_11110_10001_10001_11110;
            "C": font_data = 35'b01110_10001_10000_10000_10000_10001_01110;
            "D": font_data = 35'b11110_10001_10001_10001_10001_10001_11110;
            "E": font_data = 35'b11111_10000_10000_11110_10000_10000_11111;
            "F": font_data = 35'b11111_10000_10000_11110_10000_10000_10000;
            "G": font_data = 35'b01110_10001_10000_10111_10001_10001_01111;
            "H": font_data = 35'b10001_10001_10001_11111_10001_10001_10001;
            "I": font_data = 35'b01110_00100_00100_00100_00100_00100_01110;
            "J": font_data = 35'b00111_00010_00010_00010_00010_10010_01100;
            "K": font_data = 35'b10001_10010_10100_11000_10100_10010_10001;
            "L": font_data = 35'b10000_10000_10000_10000_10000_10000_11111;
            "M": font_data = 35'b10001_11011_10101_10101_10001_10001_10001;
            "N": font_data = 35'b10001_10001_11001_10101_10011_10001_10001;
            "O": font_data = 35'b01110_10001_10001_10001_10001_10001_01110;
            "P": font_data = 35'b11110_10001_10001_11110_10000_10000_10000;
            "Q": font_data = 35'b01110_10001_10001_10001_10101_10010_01101;
            "R": font_data = 35'b11110_10001_10001_11110_10100_10010_10001;
            "S": font_data = 35'b01111_10000_10000_01110_00001_00001_11110;
            "T": font_data = 35'b11111_00100_00100_00100_00100_00100_00100;
            "U": font_data = 35'b10001_10001_10001_10001_10001_10001_01110;
            "V": font_data = 35'b10001_10001_10001_10001_10001_01010_00100;
            "W": font_data = 35'b10001_10001_10001_10101_10101_10101_01010;
            "X": font_data = 35'b10001_10001_01010_00100_01010_10001_10001;
            "Y": font_data = 35'b10001_10001_10001_01010_00100_00100_00100;
            "Z": font_data = 35'b11111_00001_00010_00100_01000_10000_11111;
            
            // Space
            " ": font_data = 35'b00000_00000_00000_00000_00000_00000_00000;
            
            default: font_data = 35'b00000_00000_00000_00000_00000_00000_00000;
        endcase
    end

endmodule
